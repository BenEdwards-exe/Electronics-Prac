Prac4_cmos

Vdd 3 0 5
Vi 1 0 DC

MP 2 1 3 3 PMOSL
ML 2 1 0 0 NMOSD


.model PMOSL PMOS(LEVEL=1 VTO=-1.2 KP=60u)
.model NMOSD NMOS(LEVEL=1 VTO=1 KP=60u)

.DC Vi 0 5 0.05

.control
run
plot v(1), v(2)
plot i(Vdd)
.endc

.end